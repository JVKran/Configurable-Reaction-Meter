-- embedded_system_ssd_controller.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity embedded_system_ssd_controller is
	port (
		resetn     : in  std_logic                     := '0';             --    clock_reset.reset_n
		address    : in  std_logic                     := '0';             -- avalon_slave_0.address
		write      : in  std_logic                     := '0';             --               .write
		chipselect : in  std_logic                     := '0';             --               .chipselect
		writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --               .writedata
		byteenable : in  std_logic_vector(3 downto 0)  := (others => '0'); --               .byteenable
		clock      : in  std_logic                     := '0';             --     clock_sink.clk
		Q_export   : out std_logic_vector(47 downto 0)                     --    conduit_end.readdata
	);
end entity embedded_system_ssd_controller;

architecture rtl of embedded_system_ssd_controller is
	component reg32_avalon_interface is
		port (
			resetn     : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic                     := 'X';             -- address
			write      : in  std_logic                     := 'X';             -- write
			chipselect : in  std_logic                     := 'X';             -- chipselect
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clock      : in  std_logic                     := 'X';             -- clk
			Q_export   : out std_logic_vector(47 downto 0)                     -- readdata
		);
	end component reg32_avalon_interface;

begin

	ssd_controller : component reg32_avalon_interface
		port map (
			resetn     => resetn,     --    clock_reset.reset_n
			address    => address,    -- avalon_slave_0.address
			write      => write,      --               .write
			chipselect => chipselect, --               .chipselect
			writedata  => writedata,  --               .writedata
			byteenable => byteenable, --               .byteenable
			clock      => clock,      --     clock_sink.clk
			Q_export   => Q_export    --    conduit_end.readdata
		);

end architecture rtl; -- of embedded_system_ssd_controller
