-- embedded_system_response_time_meter_0.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity embedded_system_response_time_meter_0 is
	port (
		resetn   : in  std_logic                     := '0';             --         clock_reset.reset_n
		read     : in  std_logic                     := '0';             --      avalon_slave_0.read
		address  : in  std_logic                     := '0';             --                    .address
		readdata : out std_logic_vector(15 downto 0);                    --                    .readdata
		clock    : in  std_logic                     := '0';             --          clock_sink.clk
		leds     : out std_logic_vector(9 downto 0);                     --     led_conduit_end.leds_conduit
		buttons  : in  std_logic_vector(1 downto 0)  := (others => '0'); -- buttons_conduit_end.buttons_conduit
		irq      : out std_logic                                         --    interrupt_sender.irq
	);
end entity embedded_system_response_time_meter_0;

architecture rtl of embedded_system_response_time_meter_0 is
	component reg32_avalon_interface is
		port (
			resetn   : in  std_logic                     := 'X';             -- reset_n
			read     : in  std_logic                     := 'X';             -- read
			address  : in  std_logic                     := 'X';             -- address
			readdata : out std_logic_vector(15 downto 0);                    -- readdata
			clock    : in  std_logic                     := 'X';             -- clk
			leds     : out std_logic_vector(9 downto 0);                     -- leds_conduit
			buttons  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- buttons_conduit
			irq      : out std_logic                                         -- irq
		);
	end component reg32_avalon_interface;

begin

	response_time_meter_0 : component reg32_avalon_interface
		port map (
			resetn   => resetn,   --         clock_reset.reset_n
			read     => read,     --      avalon_slave_0.read
			address  => address,  --                    .address
			readdata => readdata, --                    .readdata
			clock    => clock,    --          clock_sink.clk
			leds     => leds,     --     led_conduit_end.leds_conduit
			buttons  => buttons,  -- buttons_conduit_end.buttons_conduit
			irq      => irq       --    interrupt_sender.irq
		);

end architecture rtl; -- of embedded_system_response_time_meter_0
